LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY memScor IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=130;
					ADDR_WIDTH	:	INTEGER:=5);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF memScor IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000011111111111100000000001111111110000000111111111100000011111111111111000000111111111111110000000000000000000000",
"0000000000000000000111100000011100000000011110000000000001111000011110000011111000000111100000111110000000000000000000000000000000",
"0000000000000000001111000000011111000001111100000000000001110000011110000011111000000011110000111100000000000001111000000000000000",
"0000000000000000001111000000011111000001110000000000000111100000001111100011111000000011110000111100000000000001111000000000000000",
"0000000000000000001111000000000000000111110000000000000111100000000111100011111000000011110000111100000000000001111000000000000000",
"0000000000000000001111000000000000000111110000000000000111100000000111100011111000000011110000111111111111100000000000000000000000",
"0000000000000000000111111111111100000111110000000000000111100000000111100011111000000011110000111111111111110000000000000000000000",
"0000000000000000000011111111111100000111110000000000000111100000000111100011111111111111000000111110000000000000000000000000000000",
"0000000000000000000000000000011111000111110000000000000111100000000111100011111111111111000000111100000000000000000000000000000000",
"0000000000000000000000000000011111000111110000000000000111100000000111100011111001111100000000111100000000000001111000000000000000",
"0000000000000000001111000000011111000011110000000000000111100000001111100011111000011100000000111100000000000001111000000000000000",
"0000000000000000001111000000011111000001111100000000000011110000011110000011111000001111000000111100000000000001111000000000000000",
"0000000000000000001111000000011110000001111100000000000001111000011110000011111000001111000000111100000000000001111000000000000000",
"0000000000000000000111111111111100000000001111111110000000111111111100000011111000000011110000111111111111110000000000000000000000",
"0000000000000000000011111111111100000000001111111110000000111111111000000011111000000011110000111111111111110000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

	BEGIN 

	--WRITE PROCESS
   read_process: PROCESS(clk)
	BEGIN 
		   IF (rising_edge(clk)) THEN
			data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;