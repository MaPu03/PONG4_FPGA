LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY memnum IS
	GENERIC (	DATA_WIDTH	:	INTEGER:=290;
					ADDR_WIDTH	:	INTEGER:=5);
	PORT (	clk		:	IN  STD_LOGIC;
				addr		:	IN  STD_LOGIC_VECTOR(ADDR_WIDTH-1 DOWNTO 0);
				r_data	:	OUT STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0));
END ENTITY;
-----------------------------------
ARCHITECTURE funtional OF memnum IS
----------------------------------- Build of memory
	TYPE mem_2d_type IS ARRAY (0 TO 2**ADDR_WIDTH-1) OF STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	SIGNAL ram	:	mem_2d_type;
	SIGNAL data_reg	:	STD_LOGIC_VECTOR(DATA_WIDTH-1 DOWNTO 0);
	
----------------------------------- Contents
	CONSTANT DATA_ROM: mem_2d_type:=("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000001111111111100000000000000000000011111000000000000000000011111111111111000000000000000111111111111110000000000000000000000001111100000000000011111111111111111110000000000001111111111111100000000000000111111111111111100000000000000111111111111110000000000000001111111111111100000000",
"00000000001111111111100000000000000000000111111000000000000000000011111111111111000000000000000111111111111110000000000000000000000001111100000000000011111111111111111110000000000001111111111111100000000000000111111111111111100000000000000111111111111110000000000000001111111111111100000000",
"00000000011110000011110000000000000000111111111000000000000000000011111111111111000000000000000111111111111110000000000000000000000111111100000000000011111111111111111100000000000001111111111111100000000000000111111111111111100000000000000111111111111110000000000000001111111111111100000000",
"00000000111100000011110000000000000000111111111000000000000000001111100000000111110000000000111110000000001111100000000000000000000111111100000000000011111000000000000000000000000111110000000000000000000000000000000000001111100000000000011111000000001111100000000001111100000000011111000000",
"00000000111100001111110000000000000000111111111000000000000000001111100000000111110000000000111110000000001111100000000000000000011111111100000000000011111000000000000000000000000111110000000000000000000000000000000000001111100000000000011111000000001111100000000001111110000000011111000000",
"00000011111000001100111100000000000000000011111000000000000000001111100000000111110000000000111110000000001111100000000000000000011111111100000000000011111000000000000000000000000111110000000000000000000000000000000000001111100000000000011111000000001111100000000001111110000000011111000000",
"00000011111000001100111100000000000000000011111000000000000000000000000000000111110000000000000000000000001111100000000000000000111011111100000000000011111000000000000000000000000111110000000000000000000000000000000000001111100000000000011111000000001111100000000001111110000000011111000000",
"00000011111000001100111100000000000000000011111000000000000000000000000000000111110000000000000000000000001111100000000000000011110001111100000000000000111111111111110000000000000111110000000000000000000000000000000000011100000000000000011111000000001111100000000001111110000000011111000000",
"00000011111000111000111100000000000000000011111000000000000000000000000000000111110000000000000001111111111110000000000000000011110001111100000000000000011111111111110000000000000111111111111111100000000000000000000000111100000000000000000111111111111110000000000001111100000000011111000000",
"00000011111000110000111100000000000000000011111000000000000000000011111111111111000000000000000011111111111100000000000000001111000001111100000000000000011111111111110000000000000111111111111111100000000000000000000000111100000000000000000111111111111110000000000000111110000000011111000000",
"00000011111000110000111100000000000000000011111000000000000000000011111111111111000000000000000001111111111110000000000000001111000001111100000000000000000000000000111110000000000111111111111111100000000000000000000011110000000000000000000111111111111110000000000000001111111111111111000000",
"00000011111000110000111100000000000000000011111000000000000000000011111111111111000000000000000000000000001111100000000001111100000001111100000000000000000000000000111110000000000111110000000011111100000000000000000011110000000000000000011111000000001111100000000000001111111111111111000000",
"00000011111001110000111100000000000000000011111000000000000000001111100000000000000000000000000000000000001111100000000001111100000001111100000000000000000000000000111110000000000111110000000011111100000000000000011111000000000000000000011111000000001111100000000000001111111111111111000000",
"00000011111011000000111100000000000000000011111000000000000000001111100000000000000000000000000000000000001111100000000001111110000011111100000000000011111000000000111110000000000111110000000011111100000000000000011111000000000000000000011111000000001111100000000000000000000000011111000000",
"00000011111011000000111100000000000000000011111000000000000000001111100000000000000000000000000000000000001111100000000001111111111111111111110000000011111000000000111110000000000111110000000011111100000000000000011111000000000000000000011111000000001111100000000000000000000000011111000000",
"00000011111111000011111100000000000000000011111000000000000000001111100000000000000000000000111110000000001111100000000001111111111111111111110000000011111000000000111110000000000111110000000011111100000000000000011111000000000000000000011111000000001111100000000000000000000000011111000000",
"00000000111111000011110000000000000000000011111000000000000000001111100000000000000000000000111110000000001111100000000000000000000011111100000000000011111000000000111110000000000111110000000011111100000000000000011111000000000000000000011111000000001111100000000000000000000000011111000000",
"00000000111100000011110000000000000000000011111000000000000000001111100000000000000000000000111110000000001111100000000000000000000001111100000000000011111000000000111110000000000111110000000011111100000000000000011111000000000000000000011111000000001111100000000000000000000000011111000000",
"00000000001111111111100000000000000000000111111000000000000000001111111111111111110000000000000111111111111110000000000000000000000001111100000000000000111111111111110000000000000001111111111111100000000000000000011111000000000000000000000111111111111110000000000000001111111111111100000000",
"00000000001111111111100000000000000000111111111111000000000000001111111111111111110000000000000111111111111110000000000000000000000001111100000000000000011111111111110000000000000001111111111111100000000000000000011111000000000000000000000111111111111110000000000000001111111111111100000000",
"00000000001111111111000000000000000000111111111111000000000000001111111111111111110000000000000111111111111100000000000000000000000001111100000000000000011111111111110000000000000001111111111111100000000000000000011111000000000000000000000111111111111110000000000000001111111111111100000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

	BEGIN 

	--WRITE PROCESS
   read_process: PROCESS(clk)
	BEGIN 
		   IF (rising_edge(clk)) THEN
			data_reg <= DATA_ROM(to_integer(unsigned(addr)));
		END IF;
	END PROCESS;
	--READ 
	r_data <= data_reg;
 END ARCHITECTURE funtional;